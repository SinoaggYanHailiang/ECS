library verilog;
use verilog.vl_types.all;
entity Ctr_UART is
    port(
        clk_50m         : in     vl_logic;
        rst             : in     vl_logic;
        DataRX_1        : in     vl_logic_vector(7 downto 0);
        DataRX_2        : in     vl_logic_vector(7 downto 0);
        DataRX_3        : in     vl_logic_vector(7 downto 0);
        DataRX_4        : in     vl_logic_vector(7 downto 0);
        DataRX_5        : in     vl_logic_vector(7 downto 0);
        AddrR_O         : in     vl_logic_vector(7 downto 0);
        AddrR_O_1       : in     vl_logic_vector(7 downto 0);
        Data_O_AD9244   : in     vl_logic_vector(13 downto 0);
        Data_O_AD9244_1 : in     vl_logic_vector(13 downto 0);
        Data_send_FFT   : in     vl_logic_vector(27 downto 0);
        Data_send_FFT_1 : in     vl_logic_vector(27 downto 0);
        mean_ADC1       : in     vl_logic_vector(13 downto 0);
        mean_ADC2       : in     vl_logic_vector(13 downto 0);
        flag_OverFlow_1 : in     vl_logic;
        flag_OverFlow   : in     vl_logic;
        rdy_R_AD9244    : in     vl_logic;
        rdy_R_AD9244_1  : in     vl_logic;
        rdy_W_AD9244    : in     vl_logic;
        DIO_OUT1        : out    vl_logic_vector(7 downto 0);
        DIO_OUT2        : out    vl_logic_vector(7 downto 0);
        DIO_OUT3        : out    vl_logic_vector(7 downto 0);
        Sel_WaveFunc    : out    vl_logic_vector(2 downto 0);
        DutyCyc         : out    vl_logic_vector(13 downto 0);
        freq_incr       : out    vl_logic_vector(11 downto 0);
        Amp_DAC904      : out    vl_logic_vector(15 downto 0);
        Bias_DAC904     : out    vl_logic_vector(15 downto 0);
        cnt_DAC904      : out    vl_logic_vector(39 downto 0);
        WriteEn_ADC     : out    vl_logic;
        ADCM_Length     : out    vl_logic_vector(7 downto 0);
        AddrFFT_ADC     : out    vl_logic_vector(7 downto 0);
        Flag_ReadADC_Samp: out    vl_logic;
        Flag_ReadADC_Samp_1: out    vl_logic;
        R_Restart_ADC   : out    vl_logic;
        R_Restart_ADC_1 : out    vl_logic;
        ADCR_Length     : out    vl_logic_vector(15 downto 0);
        ADCR_Length_1   : out    vl_logic_vector(15 downto 0);
        ReadFFTEn_ADC   : out    vl_logic;
        ReadFFTEn_ADC_1 : out    vl_logic;
        cnt_AD9244_W    : out    vl_logic_vector(39 downto 0);
        rst_sys         : out    vl_logic;
        DataTX_1        : out    vl_logic_vector(7 downto 0);
        DataTX_2        : out    vl_logic_vector(7 downto 0);
        DataTX_3        : out    vl_logic_vector(7 downto 0);
        DataTX_4        : out    vl_logic_vector(7 downto 0);
        EnTxData        : out    vl_logic
    );
end Ctr_UART;
