library verilog;
use verilog.vl_types.all;
entity tb_ecs is
end tb_ecs;
